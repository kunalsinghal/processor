-------------------------------------------------------
 --! @file MAUnit.vhdl
 --! @author Kunal Singhal and Swapnil Palash
 --! @brief This file for the implementation of a memory for the processor
 -------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--! This is the unit that implements a RAM. 
entity MAUnit is
	port(
		--! clk is the CLOCK coming the the unit
		clk: in std_logic;
		--! The value to stored in case of a store instruction
		op2, 
		--! aluR stores the address of the memory location to be accessed
		aluR: in std_logic_vector(31 downto 0); 
		--! a boolean signal generated by Control Unit to determine if this is a store instruction
		isSt, 
		--! a boolean signal generated by Control Unit to determine if this is a load instruction
		isLd: in boolean;
		--! output signal which contains the value stored in the memory location accessed in case of a load instruction 
		ldResult: out std_logic_vector(31 downto 0));
end entity MAUnit;

--! DM is the architecture of the Memory Unit
architecture DM of MAUnit is
	--! This is a RAM of 32768 bits that is 4096 bytes
	signal memory: std_logic_vector(32767 downto 0);
begin
	--! If there is a store instruction then this process stores the value of op2 in the required memory location
	--! If there is a load instruction then the value of required memory location is loaded into ldResult signal
	
	ldResult<=memory(to_integer(unsigned(aluR))*8+31 downto to_integer(unsigned(aluR))*8) when (isLd and (memory'event or aluR'event or isLd'event));
	
	process
	begin
		-- This line is added for the signals to get stablized
		wait until ( op2'stable(6 ns) and aluR'stable(6 ns) and isSt'stable(6 ns) and isLd'stable(6 ns));

		if (isSt and clk'event and clk='0') then 
			memory(to_integer(unsigned(aluR))*8+31 downto to_integer(unsigned(aluR))*8)<= op2;
		else null;
		end if;
	end process;
end DM;
